module array_2d_mem();
	
	reg [7:0]a[0:15][3:0];
	integer i;

	initial
		begin
		a [0] [1] [5]= 8;

			
